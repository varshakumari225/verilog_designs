module counter(input clk,rst,load,input [3:0]data,output reg [3:0]count);
  always @(posedge clk) begin
    if(rst)
      count=4'b0;
    else if (load)
      count=data;
    else
      count=count+1;
  end
endmodule
